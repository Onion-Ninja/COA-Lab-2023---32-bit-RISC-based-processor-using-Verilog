module and_gate(
    input a,
    input b,
    output wire c
);

assign c = a & b;

endmodule